** sch_path: /home/rjridle/test_current_mirror.sch
**.subckt test_current_mirror
x1 net2 current_mirror
XM1 net1 net2 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
Vdrain_current net1 GND 0
.save  i(vdrain_current)
**** begin user architecture code

.lib /import/angmar1/repos/openpdk/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt



.tran 0.1u 5u
.save all


**** end user architecture code
**.ends

* expanding   symbol:  current_mirror.sym # of pins=1
** sym_path: /home/rjridle/current_mirror.sym
** sch_path: /home/rjridle/current_mirror.sch
.subckt current_mirror  Vbias
*.opin Vbias
XM1 Vbias Vbias VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
I0 Vbias GND 3u
.ends

.GLOBAL VDD
.GLOBAL GND
.end
